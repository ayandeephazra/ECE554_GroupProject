module DM(clk,addr,re,we,wrt_data,rd_data);

/////////////////////////////////////////////////////////
// Data memory.  Single ported, can read or write but //
// not both in a single cycle.  Precharge on clock   //
// high, read/write on clock low.                   //
/////////////////////////////////////////////////////
input clk;
input [9:0] addr;
input re;				// asserted when instruction read desired
input we;				// asserted when write desired
input [16:0] wrt_data;	// data to be written

output reg [16:0] rd_data;	//output of data memory

// 2K 16-bit memory
reg [16:0]data_mem[0:1023];

// ///////////////////////////////////////////////
// // Model read, data is flopped on clock low //
// /////////////////////////////////////////////

always_ff @ (negedge clk)
  if (re && ~we)
    rd_data <= data_mem[addr];

	
// ////////////////////////////////////////////////
// // Model write, data is written on clock low //
// //////////////////////////////////////////////

always_ff @( negedge clk )
  if (we && ~re)
    data_mem[addr] <= wrt_data;
  

endmodule
